module cpu(input wire clk, reset);
//Procesador sin memoria de datos de un solo ciclo

wire s_inc, we3, wez, z, pop, push, s_stack, we4;
wire [1:0] s_inm;
wire [2:0] op_alu;
wire [5:0] opcode;

//module cd(input wire clk, reset, s_inc, we3, wez, popsignal, pushsignal, s_stack, we4,
//          input wire [1:0] s_inm,
//          input wire [2:0] op_alu, 
//          output wire z, output wire [5:0] opcode);
cd camino_datos(clk, reset, s_inc, we3, wez, pop, push, s_stack, we4,
                s_inm,
                op_alu, 
                z, opcode);

//module uc(input wire [5:0] opcode, 
//          input wire z, 
//          output reg s_inc, we3, wez, pop, push, s_stack, we4,
//          output reg [1:0] s_inm,
//          output reg [2:0] op_alu);

uc unidad_control(opcode, 
                  z, 
                  s_inc, we3, wez, pop, push, s_stack, we4,
                  s_inm,
                  op_alu);
endmodule
